// RAM

module ram #(parameter BITS=32, RAMSIZE=512, ADDR=$clog2(RAMSIZE))(
	input [BITS-1:0] dataIn,
	input read,
	input write,
	input [ADDR-1:0] address,
	input clk,
	output reg [BITS-1:0] dataOut
);

	reg [BITS-1:0] RAM [0:RAMSIZE-1];
	
	
	initial begin
		// case 1: load 
		//RAM[0] <= 'b00000_0000_0000_0000000000000000000;
		//RAM[4] <= 'b00000_0001_0000_0000000000001010101;
		//RAM[85] <= 'h0000f7f7;
		
		// case 2: load
		//RAM[0] <= 'b00000_0001_0000_0000000000000000101;
	   //RAM[4] <= 'b00000_0000_0001_0000000000000100011;
	   //RAM[40] <= 'h0000f7f7;
	
		// case 3: load imm
		//RAM[0] <= 'b00000_0001_0000_0000000000000000000;
      //RAM[4] <= 'b00001_0001_0000_0000000000001010101;
		
		// case 4: load imm
		//RAM[0] <= 'b00000_0001_0000_0000000000000000101;
      //RAM[4] <= 'b00001_0000_0001_0000000000000100011;
		
		// Store Case 1
		//RAM[0] <= 'b00000_0001_0000_0000000000001010101;
      //RAM[4] <= 'b00010_0001_0000_0000000000001011010;
		
		// Store Case 2
		//RAM[0] <= 'b00000_0001_0000_0000000000001010101;
      //RAM[4] <= 'b00010_0001_0001_0000000000001011010;
		
		// addi case 1
		//RAM[0] <= 'b00000_0001_0000_0000000000000001010;
      //RAM[4] <= 'b01011_0010_0001_1111111111111111011;
      
		// andi case 2
      //RAM[0] <= 'b00000_0001_0000_0000000000000000000;
      //RAM[4] <= 'b01011_0010_0001_0000000000000011010;
		
		// ori case 2
      //RAM[0] <= 'b00000_0001_0000_0000000000000000000;
      //RAM[4] <= 'b01011_0010_0001_0000000000000011010;
		
		// BRANCH zr case 1
		//RAM[0] <= 'b00000_0010_0000_0000000000000000000;
      //RAM[4] <= 'b10010_0010_0000_0000000000000100011;
       
		// BRANCH nz case 2
      //RAM[0] <= 'b00000_0010_0000_0000000000000000001;
      //RAM[4] <= 'b10010_0010_0001_0000000000000100011;
      
		// BRANCH pl case 3
      //RAM[0] <= 'b00000_0010_0000_0000000000000000001;
      //RAM[4] <= 'b10010_0010_0010_0000000000000100011;
       
		//BRANCH brmi case 4
      //RAM[0] <= 'b00000_0010_0000_1000000000000000001;
      //RAM[4] <= 'b10010_0010_0011_0000000000000100011;
		
		// mfhi/mflo R2
		//RAM[0] <= 'b00000_0010_0000_0000000000000000111;
		//RAM[4] <= 'b00000_0010_0000_0000000000000000000;
		
		// Jump
		//RAM[0] <= 'b00000_0001_0000_0000000000000001100;
      //RAM[4] <= 'b10011_0001_0000_0000000000000000000;

		// jump jal
	   //RAM[0] <= 'b00000_0001_0000_0000000000000001100;
      //RAM[4] <= 'b10100_0001_1111_0000000000000000001;
		
		// Input
		//RAM[0] <= 'b10101_0001_0000_0000000000000000000;
		
		// Output
      //RAM[0] <= 'b00000_0001_0000_0000000000000001111;
      //RAM[4] <= 'b10110_0001_0000_0000000000000000000;
	end

	always @ (posedge clk) begin
		if(write == 1 && read == 0) begin
			RAM[address] = dataIn;
		end
		if (read == 1 && write == 0) begin 
			dataOut = RAM[address];
		end
	end
	
endmodule
